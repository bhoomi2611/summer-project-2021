module IP(input [1:64] in, output [1:64] out);
  assign out[1] = in[58];
  assign out[2] = in[50];
  assign out[3] = in[42];
  assign out[4] = in[34];
  assign out[5] = in[26];
  assign out[6] = in[18];
  assign out[7] = in[10];
  assign out[8] = in[2];
  assign out[9] = in[60];
  assign out[10] = in[52];
  assign out[11] = in[44];
  assign out[12] = in[36];
  assign out[13] = in[28];
  assign out[14] = in[20];
  assign out[15] = in[12];
  assign out[16] = in[4];
  assign out[17] = in[62];
  assign out[18] = in[54];
  assign out[19] = in[46];
  assign out[20] = in[38];
  assign out[21] = in[30];
  assign out[22] = in[22];
  assign out[23] = in[14];
  assign out[24] = in[6];
  assign out[25] = in[64];
  assign out[26] = in[56];
  assign out[27] = in[48];
  assign out[28] = in[40];
  assign out[29] = in[32];
  assign out[30] = in[24];
  assign out[31] = in[16];
  assign out[32] = in[8];
  assign out[33] = in[57];
  assign out[34] = in[49];
  assign out[35] = in[41];
  assign out[36] = in[33];
  assign out[37] = in[25];
  assign out[38] = in[17];
  assign out[39] = in[9];
  assign out[40] = in[1];
  assign out[41] = in[59];
  assign out[42] = in[51];
  assign out[43] = in[43];
  assign out[44] = in[35];
  assign out[45] = in[27];
  assign out[46] = in[19];
  assign out[47] = in[11];
  assign out[48] = in[3];
  assign out[49] = in[61];
  assign out[50] = in[53];
  assign out[51] = in[45];
  assign out[52] = in[37];
  assign out[53] = in[29];
  assign out[54] = in[21];
  assign out[55] = in[13];
  assign out[56] = in[5];
  assign out[57] = in[63];
  assign out[58] = in[55];
  assign out[59] = in[47];
  assign out[60] = in[39];
  assign out[61] = in[31];
  assign out[62] = in[23];
  assign out[63] = in[15];
  assign out[64] = in[7];
endmodule

module IP_inv(input [1:64] in, output [1:64] out);
  assign out[1] = in[40];
  assign out[2] = in[8];
  assign out[3] = in[48];
  assign out[4] = in[16];
  assign out[5] = in[56];
  assign out[6] = in[24];
  assign out[7] = in[64];
  assign out[8] = in[32];
  assign out[9] = in[39];
  assign out[10] = in[7];
  assign out[11] = in[47];
  assign out[12] = in[15];
  assign out[13] = in[55];
  assign out[14] = in[23];
  assign out[15] = in[63];
  assign out[16] = in[31];
  assign out[17] = in[38];
  assign out[18] = in[6];
  assign out[19] = in[46];
  assign out[20] = in[14];
  assign out[21] = in[54];
  assign out[22] = in[22];
  assign out[23] = in[62];
  assign out[24] = in[30];
  assign out[25] = in[37];
  assign out[26] = in[5];
  assign out[27] = in[45];
  assign out[28] = in[13];
  assign out[29] = in[53];
  assign out[30] = in[21];
  assign out[31] = in[61];
  assign out[32] = in[29];
  assign out[33] = in[36];
  assign out[34] = in[4];
  assign out[35] = in[44];
  assign out[36] = in[12];
  assign out[37] = in[52];
  assign out[38] = in[20];
  assign out[39] = in[60];
  assign out[40] = in[28];
  assign out[41] = in[35];
  assign out[42] = in[3];
  assign out[43] = in[43];
  assign out[44] = in[11];
  assign out[45] = in[51];
  assign out[46] = in[19];
  assign out[47] = in[59];
  assign out[48] = in[27];
  assign out[49] = in[34];
  assign out[50] = in[2];
  assign out[51] = in[42];
  assign out[52] = in[10];
  assign out[53] = in[50];
  assign out[54] = in[18];
  assign out[55] = in[58];
  assign out[56] = in[26];
  assign out[57] = in[33];
  assign out[58] = in[1];
  assign out[59] = in[41];
  assign out[60] = in[9];
  assign out[61] = in[49];
  assign out[62] = in[17];
  assign out[63] = in[57];
  assign out[64] = in[25];
endmodule
module DES (input[0:63] plaintxt, input[0:55] key,output[0:63] cipher);
wire [0:63] IP_txt;
wire [0:47] Exp_right;
wire [0:47] Xor_key;
wire[0:31] S_out,permut_new,new_right;
IP ins (plaintxt, IP_txt);
// initial begin
//   #10;
//   $display("%b",IP_txt);
// end
expansion inst1(IP_txt[32:63],Exp_right);
assign Xor_key={key[0:6],key[8:14],key[16:22],key[24:30],key[32:38],key[40:46],key[48:54]}^Exp_right;
// initial begin
//   #1;
//   $display("%b",Xor_key);
// end
Sbox1 i1(Xor_key[0:5],S_out[0:3]);
// initial begin
//   #1;
//   $display("%b",S_out);
// end
Sbox2 i2(Xor_key[6:11],S_out[4:7]);
Sbox3 i3(Xor_key[12:17],S_out[8:11]);
Sbox4 i4(Xor_key[18:23],S_out[12:15]);
Sbox5 i5(Xor_key[24:29],S_out[16:19]);
Sbox6 i6(Xor_key[30:35],S_out[20:23]);
Sbox7 i7(Xor_key[36:41],S_out[24:27]);
Sbox8 i8(Xor_key[42:47],S_out[28:31]);
permute inst2(S_out,permut_new);
// initial begin
//   #1;
//   $display("%b",permut_new);
// end
//reg[0:63] IP_new;
//assign IP_new= IP_txt
assign new_right=permut_new^IP_txt[0:31];
IP_inv inst3({IP_txt[32:63],new_right},cipher);
endmodule

module Sbox1(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 14;
            S[0][1] = 4;
            S[0][2] = 13;
            S[0][3] = 1;
            S[0][4] = 2;
            S[0][5] = 15;
            S[0][6] = 11;
            S[0][7] = 8;
            S[0][8] = 3;
            S[0][9] = 10;
            S[0][10] = 6;
            S[0][11] = 12;
            S[0][12] = 5;
            S[0][13] = 9;
            S[0][14] = 0;
            S[0][15] = 7;
            S[1][0] = 0;
            S[1][1] = 15;
            S[1][2] = 7;
            S[1][3] = 4;
            S[1][4] = 14;
            S[1][5] = 2;
            S[1][6] = 13;
            S[1][7] = 1;
            S[1][8] = 10;
            S[1][9] = 6;
            S[1][10] = 12;
            S[1][11] = 11;
            S[1][12] = 9;
            S[1][13] = 5;
            S[1][14] = 3;
            S[1][15] = 8;
            S[2][0] = 4;
            S[2][1] = 1;
            S[2][2] = 14;
            S[2][3] = 8;
            S[2][4] = 13;
            S[2][5] = 6;
            S[2][6] = 2;
            S[2][7] = 11;
            S[2][8] = 15;
            S[2][9] = 12;
            S[2][10] = 9;
            S[2][11] = 7;
            S[2][12] = 3;
            S[2][13] = 10;
            S[2][14] = 5;
            S[2][15] = 0;
            S[3][0] = 15;
            S[3][1] = 12;
            S[3][2] = 8;
            S[3][3] = 2;
            S[3][4] = 4;
            S[3][5] = 9;
            S[3][6] = 1;
            S[3][7] = 7;
            S[3][8] = 5;
            S[3][9] = 11;
            S[3][10] = 3;
            S[3][11] = 14;
            S[3][12] = 10;
            S[3][13] = 0;
            S[3][14] = 6;
            S[3][15] = 13;
        
end
endmodule

module Sbox2(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 15;
            S[0][1] = 1;
            S[0][2] = 8;
            S[0][3] = 14;
            S[0][4] = 6;
            S[0][5] = 11;
            S[0][6] = 3;
            S[0][7] = 4;
            S[0][8] = 9;
            S[0][9] = 7;
            S[0][10] = 2;
            S[0][11] = 13;
            S[0][12] = 12;
            S[0][13] = 0;
            S[0][14] = 5;
            S[0][15] = 10;
            S[1][0] = 3;
            S[1][1] = 13;
            S[1][2] = 4;
            S[1][3] = 7;
            S[1][4] = 15;
            S[1][5] = 2;
            S[1][6] = 8;
            S[1][7] = 14;
            S[1][8] = 12;
            S[1][9] = 0;
            S[1][10] = 1;
            S[1][11] = 10;
            S[1][12] = 6;
            S[1][13] = 9;
            S[1][14] = 11;
            S[1][15] = 5;
            S[2][0] = 0;
            S[2][1] = 14;
            S[2][2] = 7;
            S[2][3] = 11;
            S[2][4] = 10;
            S[2][5] = 4;
            S[2][6] = 13;
            S[2][7] = 1;
            S[2][8] = 5;
            S[2][9] = 8;
            S[2][10] = 12;
            S[2][11] = 6;
            S[2][12] = 9;
            S[2][13] = 3;
            S[2][14] = 2;
            S[2][15] = 15;
            S[3][0] = 13;
            S[3][1] = 8;
            S[3][2] = 10;
            S[3][3] = 1;
            S[3][4] = 3;
            S[3][5] = 15;
            S[3][6] = 4;
            S[3][7] = 2;
            S[3][8] = 11;
            S[3][9] = 6;
            S[3][10] = 7;
            S[3][11] = 12;
            S[3][12] = 0;
            S[3][13] = 5;
            S[3][14] = 14;
            S[3][15] = 9;
 
end
endmodule

module Sbox3(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 10;
            S[0][1] = 0;
            S[0][2] = 9;
            S[0][3] = 14;
            S[0][4] = 6;
            S[0][5] = 3;
            S[0][6] = 15;
            S[0][7] = 5;
            S[0][8] = 1;
            S[0][9] = 13;
            S[0][10] = 12;
            S[0][11] = 7;
            S[0][12] = 11;
            S[0][13] = 4;
            S[0][14] = 2;
            S[0][15] = 8;
            S[1][0] = 13;
            S[1][1] = 7;
            S[1][2] = 0;
            S[1][3] = 9;
            S[1][4] = 3;
            S[1][5] = 4;
            S[1][6] = 6;
            S[1][7] = 10;
            S[1][8] = 2;
            S[1][9] = 8;
            S[1][10] = 5;
            S[1][11] = 14;
            S[1][12] = 12;
            S[1][13] = 11;
            S[1][14] = 15;
            S[1][15] = 1;
            S[2][0] = 13;
            S[2][1] = 6;
            S[2][2] = 4;
            S[2][3] = 9;
            S[2][4] = 8;
            S[2][5] = 15;
            S[2][6] = 3;
            S[2][7] = 0;
            S[2][8] = 11;
            S[2][9] = 1;
            S[2][10] = 2;
            S[2][11] = 12;
            S[2][12] = 5;
            S[2][13] = 10;
            S[2][14] = 14;
            S[2][15] = 7;
            S[3][0] = 1;
            S[3][1] = 10;
            S[3][2] = 13;
            S[3][3] = 0;
            S[3][4] = 6;
            S[3][5] = 9;
            S[3][6] = 8;
            S[3][7] = 7;
            S[3][8] = 4;
            S[3][9] = 15;
            S[3][10] = 14;
            S[3][11] = 3;
            S[3][12] = 11;
            S[3][13] = 5;
            S[3][14] = 2;
            S[3][15] = 12;

end
endmodule

module Sbox4(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 7;
            S[0][1] = 13;
            S[0][2] = 14;
            S[0][3] = 3;
            S[0][4] = 0;
            S[0][5] = 6;
            S[0][6] = 9;
            S[0][7] = 10;
            S[0][8] = 1;
            S[0][9] = 2;
            S[0][10] = 8;
            S[0][11] = 5;
            S[0][12] = 11;
            S[0][13] = 12;
            S[0][14] = 4;
            S[0][15] = 15;
            S[1][0] = 13;
            S[1][1] = 8;
            S[1][2] = 11;
            S[1][3] = 5;
            S[1][4] = 6;
            S[1][5] = 15;
            S[1][6] = 0;
            S[1][7] = 3;
            S[1][8] = 4;
            S[1][9] = 7;
            S[1][10] = 2;
            S[1][11] = 12;
            S[1][12] = 1;
            S[1][13] = 10;
            S[1][14] = 14;
            S[1][15] = 9;
            S[2][0] = 10;
            S[2][1] = 6;
            S[2][2] = 9;
            S[2][3] = 0;
            S[2][4] = 12;
            S[2][5] = 11;
            S[2][6] = 7;
            S[2][7] = 13;
            S[2][8] = 15;
            S[2][9] = 1;
            S[2][10] = 3;
            S[2][11] = 14;
            S[2][12] = 5;
            S[2][13] = 2;
            S[2][14] = 8;
            S[2][15] = 4;
            S[3][0] = 3;
            S[3][1] = 15;
            S[3][2] = 0;
            S[3][3] = 6;
            S[3][4] = 10;
            S[3][5] = 1;
            S[3][6] = 13;
            S[3][7] = 8;
            S[3][8] = 9;
            S[3][9] = 4;
            S[3][10] = 5;
            S[3][11] = 11;
            S[3][12] = 12;
            S[3][13] = 7;
            S[3][14] = 2;
            S[3][15] = 14;
end
endmodule

module Sbox5(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 2;
            S[0][1] = 12;
            S[0][2] = 4;
            S[0][3] = 1;
            S[0][4] = 7;
            S[0][5] = 10;
            S[0][6] = 11;
            S[0][7] = 6;
            S[0][8] = 8;
            S[0][9] = 5;
            S[0][10] = 3;
            S[0][11] = 15;
            S[0][12] = 13;
            S[0][13] = 0;
            S[0][14] = 14;
            S[0][15] = 9;
            S[1][0] = 14;
            S[1][1] = 11;
            S[1][2] = 2;
            S[1][3] = 12;
            S[1][4] = 4;
            S[1][5] = 7;
            S[1][6] = 13;
            S[1][7] = 1;
            S[1][8] = 5;
            S[1][9] = 0;
            S[1][10] = 15;
            S[1][11] = 10;
            S[1][12] = 3;
            S[1][13] = 9;
            S[1][14] = 8;
            S[1][15] = 6;
            S[2][0] = 4;
            S[2][1] = 2;
            S[2][2] = 1;
            S[2][3] = 11;
            S[2][4] = 10;
            S[2][5] = 13;
            S[2][6] = 7;
            S[2][7] = 8;
            S[2][8] = 15;
            S[2][9] = 9;
            S[2][10] = 12;
            S[2][11] = 5;
            S[2][12] = 6;
            S[2][13] = 3;
            S[2][14] = 0;
            S[2][15] = 14;
            S[3][0] = 11;
            S[3][1] = 8;
            S[3][2] = 12;
            S[3][3] = 7;
            S[3][4] = 1;
            S[3][5] = 14;
            S[3][6] = 2;
            S[3][7] = 13;
            S[3][8] = 6;
            S[3][9] = 15;
            S[3][10] = 0;
            S[3][11] = 9;
            S[3][12] = 10;
            S[3][13] = 4;
            S[3][14] = 5;
            S[3][15] = 3;
end
endmodule

module Sbox6(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 12;
            S[0][1] = 1;
            S[0][2] = 10;
            S[0][3] = 15;
            S[0][4] = 9;
            S[0][5] = 2;
            S[0][6] = 6;
            S[0][7] = 8;
            S[0][8] = 0;
            S[0][9] = 13;
            S[0][10] = 3;
            S[0][11] = 4;
            S[0][12] = 14;
            S[0][13] = 7;
            S[0][14] = 5;
            S[0][15] = 11;
            S[1][0] = 10;
            S[1][1] = 15;
            S[1][2] = 4;
            S[1][3] = 2;
            S[1][4] = 7;
            S[1][5] = 12;
            S[1][6] = 9;
            S[1][7] = 5;
            S[1][8] = 6;
            S[1][9] = 1;
            S[1][10] = 13;
            S[1][11] = 14;
            S[1][12] = 0;
            S[1][13] = 11;
            S[1][14] = 3;
            S[1][15] = 8;
            S[2][0] = 9;
            S[2][1] = 14;
            S[2][2] = 15;
            S[2][3] = 5;
            S[2][4] = 2;
            S[2][5] = 8;
            S[2][6] = 12;
            S[2][7] = 3;
            S[2][8] = 7;
            S[2][9] = 0;
            S[2][10] = 4;
            S[2][11] = 10;
            S[2][12] = 1;
            S[2][13] = 13;
            S[2][14] = 11;
            S[2][15] = 6;
            S[3][0] = 4;
            S[3][1] = 3;
            S[3][2] = 2;
            S[3][3] = 12;
            S[3][4] = 9;
            S[3][5] = 5;
            S[3][6] = 15;
            S[3][7] = 10;
            S[3][8] = 11;
            S[3][9] = 14;
            S[3][10] = 1;
            S[3][11] = 7;
            S[3][12] = 6;
            S[3][13] = 0;
            S[3][14] = 8;
            S[3][15] = 13;
end
endmodule

module Sbox7(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 4;
            S[0][1] = 11;
            S[0][2] = 2;
            S[0][3] = 14;
            S[0][4] = 15;
            S[0][5] = 0;
            S[0][6] = 8;
            S[0][7] = 13;
            S[0][8] = 3;
            S[0][9] = 12;
            S[0][10] = 9;
            S[0][11] = 7;
            S[0][12] = 5;
            S[0][13] = 10;
            S[0][14] = 6;
            S[0][15] = 1;
            S[1][0] = 13;
            S[1][1] = 0;
            S[1][2] = 11;
            S[1][3] = 7;
            S[1][4] = 4;
            S[1][5] = 9;
            S[1][6] = 1;
            S[1][7] = 10;
            S[1][8] = 14;
            S[1][9] = 3;
            S[1][10] = 5;
            S[1][11] = 12;
            S[1][12] = 2;
            S[1][13] = 15;
            S[1][14] = 8;
            S[1][15] = 6;
            S[2][0] = 1;
            S[2][1] = 4;
            S[2][2] = 11;
            S[2][3] = 13;
            S[2][4] = 12;
            S[2][5] = 3;
            S[2][6] = 7;
            S[2][7] = 14;
            S[2][8] = 10;
            S[2][9] = 15;
            S[2][10] = 6;
            S[2][11] = 8;
            S[2][12] = 0;
            S[2][13] = 5;
            S[2][14] = 9;
            S[2][15] = 2;
            S[3][0] = 6;
            S[3][1] = 11;
            S[3][2] = 13;
            S[3][3] = 8;
            S[3][4] = 1;
            S[3][5] = 4;
            S[3][6] = 10;
            S[3][7] = 7;
            S[3][8] = 9;
            S[3][9] = 5;
            S[3][10] = 0;
            S[3][11] = 15;
            S[3][12] = 14;
            S[3][13] = 2;
            S[3][14] = 3;
            S[3][15] = 12;
end
endmodule

module Sbox8(input[0:5] iput,output[0:3] s_out);
reg[0:3] S[0:3][0:15];
wire[0:1] row;
wire[0:3] col, s_out;
assign row = {iput[0],iput[5]};
assign col = iput[1:4];
assign  s_out = S[row][col];
initial begin
            S[0][0] = 13;
            S[0][1] = 2;
            S[0][2] = 8;
            S[0][3] = 4;
            S[0][4] = 6;
            S[0][5] = 15;
            S[0][6] = 11;
            S[0][7] = 1;
            S[0][8] = 10;
            S[0][9] = 9;
            S[0][10] = 3;
            S[0][11] = 14;
            S[0][12] = 5;
            S[0][13] = 0;
            S[0][14] = 12;
            S[0][15] = 7;
            S[1][0] = 1;
            S[1][1] = 15;
            S[1][2] = 13;
            S[1][3] = 8;
            S[1][4] = 10;
            S[1][5] = 3;
            S[1][6] = 7;
            S[1][7] = 4;
            S[1][8] = 12;
            S[1][9] = 5;
            S[1][10] = 6;
            S[1][11] = 11;
            S[1][12] = 0;
            S[1][13] = 14;
            S[1][14] = 9;
            S[1][15] = 2;
            S[2][0] = 7;
            S[2][1] = 11;
            S[2][2] = 4;
            S[2][3] = 1;
            S[2][4] = 9;
            S[2][5] = 12;
            S[2][6] = 14;
            S[2][7] = 2;
            S[2][8] = 0;
            S[2][9] = 6;
            S[2][10] = 10;
            S[2][11] = 13;
            S[2][12] = 15;
            S[2][13] = 3;
            S[2][14] = 5;
            S[2][15] = 8;
            S[3][0] = 2;
            S[3][1] = 1;
            S[3][2] = 14;
            S[3][3] = 7;
            S[3][4] = 4;
            S[3][5] = 10;
            S[3][6] = 8;
            S[3][7] = 13;
            S[3][8] = 15;
            S[3][9] = 12;
            S[3][10] = 9;
            S[3][11] = 0;
            S[3][12] = 3;
            S[3][13] = 5;
            S[3][14] = 6;
            S[3][15] = 11;
end
endmodule

module expansion(input[1:32] right,output[0:47] exp);
assign exp[0]=right[32];
assign exp[1]=right[1];
assign exp[2]=right[2];
assign exp[3]=right[3];
assign exp[4]=right[4];
assign exp[5]=right[5];
assign exp[6]=right[4];
assign exp[7]=right[5];
assign exp[8]=right[6];
assign exp[9]=right[7];
assign exp[10]=right[8];
assign exp[11]=right[9];
assign exp[12]=right[8];
assign exp[13]=right[9];
assign exp[14]=right[10];
assign exp[15]=right[11];
assign exp[16]=right[12];
assign exp[17]=right[13];
assign exp[18]=right[12];
assign exp[19]=right[13];
assign exp[20]=right[14];
assign exp[21]=right[15];
assign exp[22]=right[16];
assign exp[23]=right[17];
assign exp[24]=right[16];
assign exp[25]=right[17];
assign exp[26]=right[18];
assign exp[27]=right[19];
assign exp[28]=right[20];
assign exp[29]=right[21];
assign exp[30]=right[20];
assign exp[31]=right[21];
assign exp[32]=right[22];
assign exp[33]=right[23];
assign exp[34]=right[24];
assign exp[35]=right[25];
assign exp[36]=right[24];
assign exp[37]=right[25];
assign exp[38]=right[26];
assign exp[39]=right[27];
assign exp[40]=right[28];
assign exp[41]=right[29];
assign exp[42]=right[28];
assign exp[43]=right[29];
assign exp[44]=right[30];
assign exp[45]=right[31];
assign exp[46]=right[32];
assign exp[47]=right[1];
endmodule

module permute (input [1:32] in,output [1:32] out);
  assign out[1] = in [16];
  assign out[2] = in [7];
  assign out[3] = in [20];
  assign out[4] = in [21];
  assign out[5] = in [29];
  assign out[6] = in [12];
  assign out[7] = in [28];
  assign out[8] = in [17];
  assign out[9] = in [1];
  assign out[10] = in [15];
  assign out[11] = in [23];
  assign out[12] = in [26];
  assign out[13] = in [5];
  assign out[14] = in [18];
  assign out[15] = in [31];
  assign out[16] = in [10];
  assign out[17] = in [2];
  assign out[18] = in [8];
  assign out[19] = in [24];
  assign out[20] = in [14];
  assign out[21] = in [32];
  assign out[22] = in [27];
  assign out[23] = in [3];
  assign out[24] = in [9];
  assign out[25] = in [19];
  assign out[26] = in [13];
  assign out[27] = in [30];
  assign out[28] = in [6];
  assign out[29] = in [22];
  assign out[30] = in [11];
  assign out[31] = in [4];
  assign out[32] = in [25];
endmodule

module tb();

	reg[0:55] key;
	reg[0:63] plaintxt;
	wire[0:63] cipher;

DES inst( .plaintxt(plaintxt), .key(key),.cipher(cipher));

	initial
	begin
		plaintxt = 64'b1010101010101010101010101010101010101010101010101010101010101010;
        key = 56'b10101010101010101010101010101010101010101010101010111110;
        #10;
        $display("cipher: %b",cipher);
    plaintxt = 64'b0101011111011101111101111101010111010101110111110101110101011101;
        key = 56'b10101010101010101010101010101010101010101010101010101010;
        #10;
        $display("cipher: %b",cipher);
	end
endmodule